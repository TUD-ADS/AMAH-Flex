----------------------------------------------------------------------------------
-- Module Name: top_dummy - Behavioral
-- Project Name: -
-- Description: This top module has an empty Entity and do nothing
-- 
-- Dependencies: -
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;


entity top_dummy is

end top_dummy;

architecture Behavioral of top_dummy is


begin


end Behavioral;
